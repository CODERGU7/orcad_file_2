** Profile: "SCHEMATIC1-test"  [ D:\ae\exp2-schematic1-test.sim ] 

** Creating circuit file "exp2-schematic1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 10 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\exp2-SCHEMATIC1.net" 


.END
