** Profile: "SCHEMATIC1-f"  [ D:\ae\fullwave-schematic1-f.sim ] 

** Creating circuit file "fullwave-schematic1-f.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\fullwave-SCHEMATIC1.net" 


.END
