** Profile: "SCHEMATIC1-high "  [ D:\ae\fffffffffff-schematic1-high .sim ] 

** Creating circuit file "fffffffffff-schematic1-high .sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V2 0 5 .1 
+ LIN V_V1 0 15 5 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\fffffffffff-SCHEMATIC1.net" 


.END
