** Profile: "SCHEMATIC1-full"  [ D:\ae\full-SCHEMATIC1-full.sim ] 

** Creating circuit file "full-SCHEMATIC1-full.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\full-SCHEMATIC1.net" 


.END
